-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_0_0

-- Unique ID of L1 Trigger Menu:
-- dbf55acc-0e91-4249-aa8e-70981fc1ef36

-- Unique ID of firmware implementation:
-- 908122f9-a606-4fbc-aa7b-7864c383ad43

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.13.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i82 : std_logic;
    signal single_ext_i87 : std_logic;
    signal single_ext_i92 : std_logic;
    signal muon_shower0_i60 : std_logic;
    signal single_ett_i98 : std_logic;
    signal single_jet_i122 : std_logic;
    signal single_jet_i124 : std_logic;
    signal single_mu_i131 : std_logic;
    signal single_mu_i134 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref1_vme : std_logic;
    signal l1_bptx_beam_gas_ref1_vme : std_logic;
    signal l1_bptx_ref_and_vme : std_logic;
    signal l1_mu_shower_one_nominal : std_logic;
    signal l1_ett2000 : std_logic;
    signal l1_single_jet120er2p5 : std_logic;
    signal l1_single_jet35 : std_logic;
    signal l1_single_mu0_emtf : std_logic;
    signal l1_single_mu22_bmtf : std_logic;
    signal l1_single_mu22_emtf : std_logic;

-- ========================================================