-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_test_invmass_div_dr

-- Unique ID of L1 Trigger Menu:
-- 3c0c7341-bcb2-4f71-9732-a11cb177c360

-- Unique ID of firmware implementation:
-- 9b489ec0-fbf4-4941-985c-52e06058d80c

-- Scale set:
-- scales_2018_08_07

-- VHDL producer version
-- v2.8.0

-- ********************************************************************
-- Changed manually for muon_muon_invmass_div_dr_condition
-- ********************************************************************

-- Signal definition of pt, eta and phi for correlation conditions.
-- Insert "signal_correlation_conditions_pt_eta_phi_cos_sin_phi.vhd.j2" as often as an ObjectType at a certain Bx is used in a correlation condition.
    signal muon_pt_integer_bx_0: diff_integer_inputs_array(0 to NR_MUON_OBJECTS-1) := (others => 0);
    signal muon_pt_vector_bx_0: diff_inputs_array(0 to NR_MUON_OBJECTS-1) := (others => (others => '0'));
    signal muon_eta_integer_bx_0: diff_integer_inputs_array(0 to NR_MUON_OBJECTS-1) := (others => 0);
    signal muon_phi_integer_bx_0: diff_integer_inputs_array(0 to NR_MUON_OBJECTS-1) := (others => 0);
    signal muon_cos_phi_bx_0: sin_cos_integer_array(0 to NR_MUON_OBJECTS-1) := (others => 0);
    signal muon_sin_phi_bx_0: sin_cos_integer_array(0 to NR_MUON_OBJECTS-1) := (others => 0);
    signal muon_eta_conv_2_muon_eta_integer_bx_0: diff_integer_inputs_array(0 to NR_MUON_OBJECTS-1) := (others => 0);
    signal muon_phi_conv_2_muon_phi_integer_bx_0: diff_integer_inputs_array(0 to NR_MUON_OBJECTS-1) := (others => 0);

-- Signal definition of differences for correlation conditions.
-- Insert "signal_correlation_conditions_differences.vhd.j2" once for correlation conditions of different ObjectTypes and Bx combinations.
    signal muon_muon_bx_0_bx_0_diff_eta_integer: dim2_max_eta_range_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => 0));
    signal muon_muon_bx_0_bx_0_diff_eta_integer_lut: diff_2dim_integer_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => 0));
    signal muon_muon_bx_0_bx_0_diff_eta_vector: deta_dphi_vector_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => (others => '0')));
    signal muon_muon_bx_0_bx_0_diff_phi_integer: dim2_max_phi_range_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => 0));
    signal muon_muon_bx_0_bx_0_diff_phi_integer_lut: diff_2dim_integer_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => 0));
    signal muon_muon_bx_0_bx_0_diff_phi_vector: deta_dphi_vector_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => (others => '0')));
    signal muon_muon_bx_0_bx_0_cosh_deta_integer : diff_2dim_integer_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => 0));
    signal muon_muon_bx_0_bx_0_cosh_deta_vector : muon_cosh_cos_vector_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => (others => '0')));
    signal muon_muon_bx_0_bx_0_cos_dphi_integer : diff_2dim_integer_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => 0));
    signal muon_muon_bx_0_bx_0_cos_dphi_vector : muon_cosh_cos_vector_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => (others => '0')));

    signal muon_muon_bx_0_bx_0_deta_bin_vector : muon_deta_bin_vector_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => (others => '0')));
    signal muon_muon_bx_0_bx_0_dphi_bin_vector : muon_dphi_bin_vector_array(0 to NR_MUON_OBJECTS-1, 0 to NR_MUON_OBJECTS-1) := (others => (others => (others => '0')));
    
-- Signal definition for muon charge correlations.
-- Insert "signal_muon_charge_correlations.vhd.j2" only once for a certain Bx combination,
-- if there is at least one muon condition or one muon-muon correlation condition.

-- Signal definition for conditions names
    signal invariant_mass_i0 : std_logic;

-- Signal definition for algorithms names
    signal l1_muon_invmass_div_dr : std_logic;

-- ========================================================
