-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_utm_0_11_test

-- Unique ID of L1 Trigger Menu:
-- 36a2b4c9-da1a-4698-be00-93a32f4e85dc

-- Unique ID of firmware implementation:
-- d6d7d469-f972-4239-8cb5-0fb4c6b13751

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.0

-- tmEventSetup version
-- v0.11.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal muon_shower2_i5 : std_logic;
    signal zdc_plus_i6 : std_logic;

-- Signal definition for algorithms names
    signal l1_zdc_plus_128 : std_logic;
    signal l1_single_mu_shower_two_loose : std_logic;

-- ========================================================