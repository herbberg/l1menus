-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_Cicada_Topo_test_v4

-- Unique ID of L1 Trigger Menu:
-- e50b8093-a248-4fd5-baf6-5b197178654a

-- Unique ID of firmware implementation:
-- 77aeb023-0ba8-4f76-920d-188621641271

-- Scale set:
-- scales_2023_12_14

-- VHDL producer version
-- v2.17.0

-- tmEventSetup version
-- v0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal cicada_trigger_i0 : std_logic;
    signal cicada_trigger_i1 : std_logic;
    signal cicada_trigger_i2 : std_logic;
    signal cicada_trigger_i3 : std_logic;
    signal cicada_trigger_i4 : std_logic;
    signal single_eg_i7 : std_logic;

-- Signal definition for algorithms names
    signal l1_cicada_4p273_and_3p0 : std_logic;
    signal l1_cicada_5p273 : std_logic;
    signal l1_cicada_142p273 : std_logic;
    signal l1_cicada_10p023 : std_logic;
    signal l1_single_eg8er2p5 : std_logic;

-- ========================================================