    signal dout : std_logic_vector(25 downto 0) := (others => '0');
    signal addr_lsb : std_logic_vector(11 DOWNTO 0) := (others => '0');

-- Signal definition for algorithms names
    signal l1_dummy : std_logic := '0';

-- ========================================================
