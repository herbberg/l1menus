-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_test_compare_gtl_struct_v6

-- Unique ID of L1 Trigger Menu:
-- fbf199b0-440e-4a10-9b8b-d4847a9b443d

-- Unique ID of firmware implementation:
-- 472e5ea1-1a83-4a99-b8d1-d66a95206ce1

-- Scale set:
-- scales_2018_08_07

-- VHDL producer version
-- v2.7.2

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
          0, -- module_index: 0, name: L1_Test_DoubleJet30_Tbpt60
          2, -- module_index: 1, name: L1_Test_DoubleJet30_Tau45_Deta_ignore_Tbpt60_OrmDr0p2
    others => 0
);

-- ========================================================