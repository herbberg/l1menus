-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_Axol1tl_Cicada_Topo_model_cut_test_v4

-- Unique ID of L1 Trigger Menu:
-- 6eae7c81-757b-45f7-878c-0ab2c2f2bdd2

-- Unique ID of firmware implementation:
-- 09c0303c-3d78-4fd5-89d5-a7426d7c7be4

-- Scale set:
-- scales_2024_01_04

-- VHDL producer version
-- v2.17.0

-- tmEventSetup version
-- v0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal cicada_trigger_i0 : std_logic;
    signal cicada_trigger_i1 : std_logic;
    signal cicada_trigger_i4 : std_logic;
    signal cicada_trigger_i6 : std_logic;

-- Signal definition for algorithms names
    signal l1_cicada_4p273_and_3p0 : std_logic;
    signal l1_cicada_10p023 : std_logic;
    signal l1_cicada_45p801 : std_logic;

-- ========================================================