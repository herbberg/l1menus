-- ========================================================
-- from VHDL producer:

-- Module ID: 2

-- Name of L1 Trigger Menu:
-- L1Menu_test_all_condition_types_v5

-- Unique ID of L1 Trigger Menu:
-- 9b8f1705-dedd-4cba-b11d-409cb9fe35e1

-- Unique ID of firmware implementation:
-- fc7bc2f8-5838-4df5-ba33-ab67aab96ba2

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.11.0

-- tmEventSetup version
-- v0.8.1

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
         54, -- module_index: 0, name: L1_DoubleMu0er2p0_SQ_OS_dR_Max1p4
        199, -- module_index: 1, name: L1_IsoEG32er2p5_Mt48
        143, -- module_index: 2, name: L1_DoubleMu3_dR_Max1p6_Jet90er2p5_dR_Max0p8
          9, -- module_index: 3, name: L1_DoubleMU20_30_MASSDR_min_10
    others => 0
);

-- ========================================================