-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_1_0_utm_0_11

-- Unique ID of L1 Trigger Menu:
-- 4539b19c-42d9-43bf-b18a-d5e88a271ad2

-- Unique ID of firmware implementation:
-- 8573c090-c2e3-4197-a299-04818e4251d0

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.0

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i1 : std_logic;
    signal single_ext_i11 : std_logic;
    signal single_ext_i6 : std_logic;
    signal muon_shower1_i15 : std_logic;
    signal single_ett_i20 : std_logic;
    signal single_jet_i60 : std_logic;
    signal single_jet_i62 : std_logic;
    signal single_mu_i70 : std_logic;
    signal single_mu_i73 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref1_vme : std_logic;
    signal l1_bptx_beam_gas_ref1_vme : std_logic;
    signal l1_bptx_ref_and_vme : std_logic;
    signal l1_mu_shower_one_tight : std_logic;
    signal l1_ett2000 : std_logic;
    signal l1_single_jet120er2p5 : std_logic;
    signal l1_single_jet35 : std_logic;
    signal l1_single_mu0_emtf : std_logic;
    signal l1_single_mu22_bmtf : std_logic;
    signal l1_single_mu22_emtf : std_logic;

-- ========================================================