-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_Axol1tl_Cicada_Topo_model_cut_test_v7

-- Unique ID of L1 Trigger Menu:
-- 5a1c2a44-d0d5-4a3b-ba17-e4223a7798bb

-- Unique ID of firmware implementation:
-- 7725cb3d-b7b8-4e1a-84e4-5280b005245f

-- Scale set:
-- scales_2024_01_04

-- VHDL producer version
-- v2.17.0

-- tmEventSetup version
-- v0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal cicada_trigger_i4 : std_logic;
    signal cicada_trigger_i6 : std_logic;
    signal topological_trigger_i11 : std_logic;

-- Signal definition for algorithms names
    signal l1_cicada_10p023 : std_logic;
    signal l1_topo_300_hh_had_v1 : std_logic;
    signal l1_cicada_45p801 : std_logic;

-- ========================================================