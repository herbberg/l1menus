-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_Cicada_Topo_test

-- Unique ID of L1 Trigger Menu:
-- e50b8093-a248-4fd5-baf6-5b197178654a

-- Unique ID of firmware implementation:
-- 5e376639-dc6d-42ec-bc44-fc07141566e4

-- Scale set:
-- scales_2023_12_14

-- VHDL producer version
-- v2.17.0

-- tmEventSetup version
-- v0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal cicada_trigger_i2 : std_logic;
    signal cicada_trigger_i4 : std_logic;

-- Signal definition for algorithms names
    signal l1_cicada_5p273 : std_logic;
    signal l1_cicada_10p023 : std_logic;

-- ========================================================