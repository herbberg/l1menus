-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_test_all_condition_types_v3

-- Unique ID of L1 Trigger Menu:
-- ad621df6-97ab-423f-baf3-0bddfb83d618

-- Unique ID of firmware implementation:
-- 42d1de01-2dd9-4e11-9083-de83a1bdad02

-- Scale set:
-- scales_2020_10_04

-- VHDL producer version
-- v2.11.0

-- tmEventSetup version
-- v0.8.1

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        410, -- module_index: 0, name: L1_ETT1200
        400, -- module_index: 1, name: L1_HTT200er
        160, -- module_index: 2, name: L1_SingleEG10er2p5
         18, -- module_index: 3, name: L1_SingleMu20
         99, -- module_index: 4, name: L1_Mu20_EG10er2p5
        194, -- module_index: 5, name: L1_SingleIsoEG32er2p5
        331, -- module_index: 6, name: L1_SingleJet12erHE
        314, -- module_index: 7, name: L1_SingleJet200
        310, -- module_index: 8, name: L1_SingleJet60
        318, -- module_index: 9, name: L1_SingleJet90er2p5
          2, -- module_index: 10, name: L1_Eg20_Jet40_ORMDR_min_2p4
        206, -- module_index: 11, name: L1_DoubleEG_20_10_er2p5
        208, -- module_index: 12, name: L1_DoubleEG_25_12_er2p5
        212, -- module_index: 13, name: L1_DoubleEG_LooseIso20_10_er2p5
        215, -- module_index: 14, name: L1_DoubleEG_LooseIso25_12_er2p5
        271, -- module_index: 15, name: L1_DoubleIsoTau32er2p1
        341, -- module_index: 16, name: L1_DoubleJet100er2p5
        218, -- module_index: 17, name: L1_DoubleLooseIsoEG24er2p1
        327, -- module_index: 18, name: L1_SingleJet120_FWD3p0
        228, -- module_index: 19, name: L1_TripleEG16er2p5
        227, -- module_index: 20, name: L1_TripleEG_18_18_12_er2p5
        305, -- module_index: 21, name: L1_Mu0upt100
        154, -- module_index: 22, name: L1_Mu0upt20ip1
        304, -- module_index: 23, name: L1_Mu0upt50
         14, -- module_index: 24, name: L1_SingleMu12_DQ_OMTF
         32, -- module_index: 25, name: L1_SingleMu16er1p5
         20, -- module_index: 26, name: L1_SingleMu22_BMTF
         25, -- module_index: 27, name: L1_SingleMu6er1p5
         27, -- module_index: 28, name: L1_SingleMu8er1p5
        307, -- module_index: 29, name: L1_SingleMuOpenupt20
        119, -- module_index: 30, name: L1_Mu3_Jet30er2p5
         40, -- module_index: 31, name: L1_DoubleMu0
         42, -- module_index: 32, name: L1_DoubleMu0_SQ_OS
         56, -- module_index: 33, name: L1_DoubleMu0er1p5_SQ_OS
         60, -- module_index: 34, name: L1_DoubleMu4_SQ_OS
         64, -- module_index: 35, name: L1_DoubleMu4p5er2p0_SQ_OS
         45, -- module_index: 36, name: L1_DoubleMu9_SQ
         47, -- module_index: 37, name: L1_DoubleMu_15_5_SQ
         49, -- module_index: 38, name: L1_DoubleMu_15_7_SQ
         72, -- module_index: 39, name: L1_TripleMu0
         73, -- module_index: 40, name: L1_TripleMu0_SQ
         75, -- module_index: 41, name: L1_TripleMu3_SQ
         78, -- module_index: 42, name: L1_TripleMu_5_3_3
         79, -- module_index: 43, name: L1_TripleMu_5_3_3_SQ
         77, -- module_index: 44, name: L1_TripleMu_5_3p5_2p5
         84, -- module_index: 45, name: L1_TripleMu_5_4_2p5_DoubleMu_5_2p5_OS_Mass_5to17
         83, -- module_index: 46, name: L1_TripleMu_5_3p5_2p5_DoubleMu_5_2p5_OS_Mass_5to17
         58, -- module_index: 47, name: L1_DoubleMu0er1p5_SQ_OS_dR_Max1p4
         61, -- module_index: 48, name: L1_DoubleMu4_SQ_OS_dR_Max1p2
        199, -- module_index: 49, name: L1_IsoEG32er2p5_Mt48
        382, -- module_index: 50, name: L1_QuadJet60er2p5
        276, -- module_index: 51, name: L1_DoubleIsoTau30er2p1_Mass_Max90
        351, -- module_index: 52, name: L1_DoubleJet30er2p5_Mass_Min300_dEta_Max1p5
        234, -- module_index: 53, name: L1_LooseIsoEG26er2p1_Jet34er2p5_dR_Min0p3
        126, -- module_index: 54, name: L1_Mu3_Jet120er2p5_dR_Max0p4
        136, -- module_index: 55, name: L1_Mu12er2p3_Jet40er2p1_dR_Max0p4_DoubleJet40er2p1_dEta_Max1p6
          0, -- module_index: 56, name: L1_DoubleJet20_30_slice_0_5_MASSDR_min_10
    others => 0
);

-- ========================================================