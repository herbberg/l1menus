-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2020_v0_1_2_with_JET_DISP_LLP_v2

-- Unique ID of L1 Trigger Menu:
-- 583970d6-daf2-445f-909e-cc79eaaf846c

-- Unique ID of firmware implementation:
-- 6b89c3ff-74a3-4b78-8cc1-dbf1cb5f2a11

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.12.0

-- tmEventSetup version
-- v0.10.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        491, -- module_index: 0, name: L1_BPTX_BeamGas_B1_VME
        483, -- module_index: 1, name: L1_BPTX_OR_Ref3_VME
        479, -- module_index: 2, name: L1_FirstCollisionInTrain
        503, -- module_index: 3, name: L1_TOTEM_1
        469, -- module_index: 4, name: L1_UnpairedBunchBptxMinus
        426, -- module_index: 5, name: L1_ETMHF150
        399, -- module_index: 6, name: L1_HTT160er
        406, -- module_index: 7, name: L1_HTT450er
         18, -- module_index: 8, name: L1_SingleMu20
         99, -- module_index: 9, name: L1_Mu20_EG10er2p5
        160, -- module_index: 10, name: L1_SingleEG10er2p5
        313, -- module_index: 11, name: L1_SingleJet180
        310, -- module_index: 12, name: L1_SingleJet60
        302, -- module_index: 13, name: L1_Mu0upt10
        301, -- module_index: 14, name: L1_Mu0upt5
        157, -- module_index: 15, name: L1_Mu0upt20ip03
        156, -- module_index: 16, name: L1_Mu0upt20ip3
        308, -- module_index: 17, name: L1_SingleMuOpenupt100
         29, -- module_index: 18, name: L1_SingleMu10er1p5
         32, -- module_index: 19, name: L1_SingleMu16er1p5
         26, -- module_index: 20, name: L1_SingleMu7er1p5
         39, -- module_index: 21, name: L1_DoubleMu0_OQ
         46, -- module_index: 22, name: L1_DoubleMu_12_5
         49, -- module_index: 23, name: L1_DoubleMu_15_7_SQ
         62, -- module_index: 24, name: L1_DoubleMu4p5_SQ_OS
        166, -- module_index: 25, name: L1_SingleEG28er1p5
        167, -- module_index: 26, name: L1_SingleEG34er2p5
        170, -- module_index: 27, name: L1_SingleEG40er2p5
        159, -- module_index: 28, name: L1_SingleEG8er2p5
        322, -- module_index: 29, name: L1_SingleJet180er2p5
          3, -- module_index: 30, name: L1_SingleMuCosmics_EMTF
        265, -- module_index: 31, name: L1_SingleTau130er2p1
         15, -- module_index: 32, name: L1_SingleMu12_DQ_EMTF
         21, -- module_index: 33, name: L1_SingleMu22_OMTF
        187, -- module_index: 34, name: L1_SingleIsoEG26er1p5
        191, -- module_index: 35, name: L1_SingleIsoEG28er1p5
        193, -- module_index: 36, name: L1_SingleIsoEG30er2p1
        194, -- module_index: 37, name: L1_SingleIsoEG32er2p5
        175, -- module_index: 38, name: L1_SingleLooseIsoEG26er2p5
        178, -- module_index: 39, name: L1_SingleLooseIsoEG28er2p5
        181, -- module_index: 40, name: L1_SingleLooseIsoEG30er2p5
        198, -- module_index: 41, name: L1_IsoEG32er2p5_Mt44
         71, -- module_index: 42, name: L1_TripleMu0_OQ
         74, -- module_index: 43, name: L1_TripleMu3
         78, -- module_index: 44, name: L1_TripleMu_5_3_3
         77, -- module_index: 45, name: L1_TripleMu_5_3p5_2p5
         83, -- module_index: 46, name: L1_TripleMu_5_3p5_2p5_DoubleMu_5_2p5_OS_Mass_5to17
         84, -- module_index: 47, name: L1_TripleMu_5_4_2p5_DoubleMu_5_2p5_OS_Mass_5to17
         89, -- module_index: 48, name: L1_QuadMu0
         90, -- module_index: 49, name: L1_QuadMu0_SQ
        205, -- module_index: 50, name: L1_DoubleEG_15_10_er2p5
        206, -- module_index: 51, name: L1_DoubleEG_20_10_er2p5
        208, -- module_index: 52, name: L1_DoubleEG_25_12_er2p5
        210, -- module_index: 53, name: L1_DoubleEG_27_14_er2p5
        342, -- module_index: 54, name: L1_DoubleJet120er2p5
        267, -- module_index: 55, name: L1_DoubleTau70er2p1
        327, -- module_index: 56, name: L1_SingleJet120_FWD3p0
        326, -- module_index: 57, name: L1_SingleJet90_FWD3p0
        214, -- module_index: 58, name: L1_DoubleEG_LooseIso22_12_er2p5
        269, -- module_index: 59, name: L1_DoubleIsoTau28er2p1
        271, -- module_index: 60, name: L1_DoubleIsoTau32er2p1
        273, -- module_index: 61, name: L1_DoubleIsoTau36er2p1
        218, -- module_index: 62, name: L1_DoubleLooseIsoEG24er2p1
        177, -- module_index: 63, name: L1_SingleLooseIsoEG28_FWD2p5
        224, -- module_index: 64, name: L1_TripleEG_16_12_8_er2p5
        226, -- module_index: 65, name: L1_TripleEG_18_17_8_er2p5
        374, -- module_index: 66, name: L1_TripleJet_105_85_75_DoubleJet_85_75_er2p5
        298, -- module_index: 67, name: L1_QuadJet36er2p5_IsoTau52er2p1
        346, -- module_index: 68, name: L1_DoubleJet112er2p3_dEta_Max1p6
         54, -- module_index: 69, name: L1_DoubleMu0er2p0_SQ_OS_dR_Max1p4
         50, -- module_index: 70, name: L1_DoubleMu_15_7_Mass_Min1
         82, -- module_index: 71, name: L1_TripleMu_5_3p5_2p5_OQ_DoubleMu_5_2p5_OQ_OS_Mass_5to17
        125, -- module_index: 72, name: L1_Mu3_Jet120er2p5_dR_Max0p8
        134, -- module_index: 73, name: L1_Mu10er2p3_Jet32er2p3_dR_Max0p4_DoubleJet32er2p3_dEta_Max1p6
        142, -- module_index: 74, name: L1_DoubleMu0_dR_Max1p6_Jet90er2p5_dR_Max0p8
        356, -- module_index: 75, name: L1_DoubleJet_100_30_DoubleJet30_Mass_Min620
        355, -- module_index: 76, name: L1_DoubleJet_90_30_DoubleJet30_Mass_Min620
        348, -- module_index: 77, name: L1_DoubleJet30er2p5_Mass_Min150_dEta_Max1p5
        350, -- module_index: 78, name: L1_DoubleJet30er2p5_Mass_Min250_dEta_Max1p5
        352, -- module_index: 79, name: L1_DoubleJet30er2p5_Mass_Min330_dEta_Max1p5
        236, -- module_index: 80, name: L1_LooseIsoEG30er2p1_Jet34er2p5_dR_Min0p3
    others => 0
);

-- ========================================================