-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2018_v4_2_0_new_scale

-- Unique ID of L1 Trigger Menu:
-- 786b195b-7fe4-4c23-a571-ac5068c6fa09

-- Unique ID of firmware implementation:
-- 16aa0ff4-bb99-4e7c-93a6-91d053a5e21c

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.12.1

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.
    signal eg_bx_0_pt_vector: diff_inputs_array(0 to NR_EG_OBJECTS-1) := (others => (others => '0'));
    signal eg_bx_0_eta_integer: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal eg_bx_0_phi_integer: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal eg_bx_0_cos_phi: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal eg_bx_0_sin_phi: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal eg_bx_0_conv_cos_phi: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal eg_bx_0_conv_sin_phi: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal eg_bx_0_eta_conv_2_muon_eta_integer: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal eg_bx_0_phi_conv_2_muon_phi_integer: integer_array(0 to NR_EG_OBJECTS-1) := (others => 0);
    signal jet_bx_0_pt_vector: diff_inputs_array(0 to NR_JET_OBJECTS-1) := (others => (others => '0'));
    signal jet_bx_0_eta_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_phi_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_cos_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_sin_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_conv_cos_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_conv_sin_phi: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_eta_conv_2_muon_eta_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal jet_bx_0_phi_conv_2_muon_phi_integer: integer_array(0 to NR_JET_OBJECTS-1) := (others => 0);
    signal mu_bx_0_pt_vector: diff_inputs_array(0 to NR_MU_OBJECTS-1) := (others => (others => '0'));
    signal mu_bx_0_upt_vector: diff_inputs_array(0 to NR_MU_OBJECTS-1) := (others => (others => '0'));
    signal mu_bx_0_eta_integer: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_phi_integer: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_eta_integer_half_res: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_phi_integer_half_res: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_cos_phi: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);
    signal mu_bx_0_sin_phi: integer_array(0 to NR_MU_OBJECTS-1) := (others => 0);

-- Signal definition for cuts of correlation conditions.
    signal eg_jet_bx_0_bx_0_deta_integer: dim2_max_eta_range_array(0 to NR_EG_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => 0));
    signal eg_jet_bx_0_bx_0_deta: deta_dphi_vector_array(0 to NR_EG_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => (others => '0')));
    signal eg_jet_bx_0_bx_0_dphi_integer: dim2_max_phi_range_array(0 to NR_EG_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => 0));
    signal eg_jet_bx_0_bx_0_dphi: deta_dphi_vector_array(0 to NR_EG_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_deta_integer: dim2_max_eta_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal mu_mu_bx_0_bx_0_deta: deta_dphi_vector_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_dphi_integer: dim2_max_phi_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal mu_mu_bx_0_bx_0_dphi: deta_dphi_vector_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_deta_integer_half_res: dim2_max_eta_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal mu_mu_bx_0_bx_0_dphi_integer_half_res: dim2_max_phi_range_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => 0));
    signal eg_jet_bx_0_bx_0_dr : dr_dim2_array(0 to NR_EG_OBJECTS-1, 0 to NR_JET_OBJECTS-1) := (others => (others => (others => '0')));
    signal mu_mu_bx_0_bx_0_dr : dr_dim2_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1) := (others => (others => (others => '0')));

-- Signal definition for muon charge correlations.
    signal ls_charcorr_double_bx_0_bx_0, os_charcorr_double_bx_0_bx_0 : std_logic_2dim_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1);
    signal ls_charcorr_triple_bx_0_bx_0, os_charcorr_triple_bx_0_bx_0 : std_logic_3dim_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1);
    signal ls_charcorr_quad_bx_0_bx_0, os_charcorr_quad_bx_0_bx_0 : std_logic_4dim_array(0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1, 0 to NR_MU_OBJECTS-1);

-- Signal definition for conditions names
    signal single_asymet_i172 : std_logic;
    signal single_asymet_i173 : std_logic;
    signal single_asymet_i174 : std_logic;
    signal single_asymet_i175 : std_logic;
    signal single_asymet_i176 : std_logic;
    signal single_asymet_i178 : std_logic;
    signal single_asymet_i179 : std_logic;
    signal single_cent0_i81 : std_logic;
    signal single_cent1_i82 : std_logic;
    signal single_cent2_i83 : std_logic;
    signal single_cent3_i84 : std_logic;
    signal single_cent4_i85 : std_logic;
    signal single_cent5_i98 : std_logic;
    signal single_cent6_i119 : std_logic;
    signal single_ext_i12 : std_logic;
    signal single_ext_i198 : std_logic;
    signal single_ext_i199 : std_logic;
    signal single_ext_i200 : std_logic;
    signal single_ext_i57 : std_logic;
    signal single_ext_i58 : std_logic;
    signal single_ext_i60 : std_logic;
    signal single_ext_i61 : std_logic;
    signal single_ext_i62 : std_logic;
    signal single_ext_i65 : std_logic;
    signal single_ext_i70 : std_logic;
    signal single_ext_i71 : std_logic;
    signal single_ext_i72 : std_logic;
    signal single_ext_i73 : std_logic;
    signal single_ext_i74 : std_logic;
    signal single_ext_i75 : std_logic;
    signal single_ext_i76 : std_logic;
    signal single_ext_i77 : std_logic;
    signal single_ext_i80 : std_logic;
    signal single_mbt0_hfm_i64 : std_logic;
    signal single_mbt1_hfm_i22 : std_logic;
    signal single_mbt0_hfp_i63 : std_logic;
    signal single_mbt1_hfp_i21 : std_logic;
    signal single_ett_i177 : std_logic;
    signal single_ett_i180 : std_logic;
    signal single_ett_i181 : std_logic;
    signal single_ett_i182 : std_logic;
    signal single_ett_i183 : std_logic;
    signal single_ett_i184 : std_logic;
    signal single_ett_i185 : std_logic;
    signal single_ett_i186 : std_logic;
    signal single_ett_i187 : std_logic;
    signal single_ett_i188 : std_logic;
    signal single_ett_i189 : std_logic;
    signal single_ett_i190 : std_logic;
    signal single_ett_i191 : std_logic;
    signal single_ett_i192 : std_logic;
    signal single_ett_i193 : std_logic;
    signal single_ett_i194 : std_logic;
    signal single_ett_i195 : std_logic;
    signal single_ett_i196 : std_logic;
    signal single_ett_i54 : std_logic;
    signal single_ett_i97 : std_logic;
    signal calo_calo_correlation_i157 : std_logic;
    signal calo_calo_correlation_i158 : std_logic;
    signal calo_calo_correlation_i159 : std_logic;
    signal calo_calo_correlation_i160 : std_logic;
    signal calo_calo_correlation_i161 : std_logic;
    signal calo_calo_correlation_i162 : std_logic;
    signal calo_calo_correlation_i163 : std_logic;
    signal calo_calo_correlation_i164 : std_logic;
    signal calo_calo_correlation_i166 : std_logic;
    signal calo_calo_correlation_i167 : std_logic;
    signal calo_calo_correlation_i168 : std_logic;
    signal calo_calo_correlation_i169 : std_logic;
    signal muon_muon_correlation_i116 : std_logic;
    signal muon_muon_correlation_i117 : std_logic;
    signal muon_muon_correlation_i118 : std_logic;
    signal double_eg_i170 : std_logic;
    signal double_eg_i171 : std_logic;
    signal double_eg_i33 : std_logic;
    signal double_eg_i34 : std_logic;
    signal double_jet_i146 : std_logic;
    signal double_jet_i147 : std_logic;
    signal double_jet_i148 : std_logic;
    signal double_jet_i149 : std_logic;
    signal double_jet_i150 : std_logic;
    signal double_mu_i113 : std_logic;
    signal double_mu_i114 : std_logic;
    signal double_mu_i115 : std_logic;
    signal double_mu_i20 : std_logic;
    signal double_mu_i23 : std_logic;
    signal single_eg_i107 : std_logic;
    signal single_eg_i108 : std_logic;
    signal single_eg_i109 : std_logic;
    signal single_eg_i110 : std_logic;
    signal single_eg_i111 : std_logic;
    signal single_eg_i112 : std_logic;
    signal single_eg_i151 : std_logic;
    signal single_eg_i152 : std_logic;
    signal single_eg_i153 : std_logic;
    signal single_eg_i154 : std_logic;
    signal single_eg_i155 : std_logic;
    signal single_eg_i156 : std_logic;
    signal single_eg_i26 : std_logic;
    signal single_eg_i27 : std_logic;
    signal single_jet_i101 : std_logic;
    signal single_jet_i102 : std_logic;
    signal single_jet_i103 : std_logic;
    signal single_jet_i104 : std_logic;
    signal single_jet_i105 : std_logic;
    signal single_jet_i106 : std_logic;
    signal single_jet_i120 : std_logic;
    signal single_jet_i121 : std_logic;
    signal single_jet_i122 : std_logic;
    signal single_jet_i123 : std_logic;
    signal single_jet_i124 : std_logic;
    signal single_jet_i125 : std_logic;
    signal single_jet_i126 : std_logic;
    signal single_jet_i127 : std_logic;
    signal single_jet_i128 : std_logic;
    signal single_jet_i129 : std_logic;
    signal single_jet_i130 : std_logic;
    signal single_jet_i131 : std_logic;
    signal single_jet_i132 : std_logic;
    signal single_jet_i133 : std_logic;
    signal single_jet_i134 : std_logic;
    signal single_jet_i135 : std_logic;
    signal single_jet_i136 : std_logic;
    signal single_jet_i137 : std_logic;
    signal single_jet_i138 : std_logic;
    signal single_jet_i139 : std_logic;
    signal single_jet_i140 : std_logic;
    signal single_jet_i141 : std_logic;
    signal single_jet_i142 : std_logic;
    signal single_jet_i143 : std_logic;
    signal single_jet_i144 : std_logic;
    signal single_jet_i145 : std_logic;
    signal single_jet_i165 : std_logic;
    signal single_jet_i35 : std_logic;
    signal single_jet_i37 : std_logic;
    signal single_mu_i10 : std_logic;
    signal single_mu_i100 : std_logic;
    signal single_mu_i11 : std_logic;
    signal single_mu_i13 : std_logic;
    signal single_mu_i14 : std_logic;
    signal single_mu_i15 : std_logic;
    signal single_mu_i4 : std_logic;
    signal single_mu_i6 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_mu_open : std_logic;
    signal l1_single_mu0 : std_logic;
    signal l1_single_mu3 : std_logic;
    signal l1_single_mu3_open_bptx_and : std_logic;
    signal l1_single_mu5 : std_logic;
    signal l1_single_mu7 : std_logic;
    signal l1_single_mu12 : std_logic;
    signal l1_double_mu_open_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_mu0 : std_logic;
    signal l1_single_eg3 : std_logic;
    signal l1_single_eg5 : std_logic;
    signal l1_double_eg2 : std_logic;
    signal l1_double_eg5 : std_logic;
    signal l1_single_jet8 : std_logic;
    signal l1_single_jet60 : std_logic;
    signal l1_ett5 : std_logic;
    signal l1_totem_1 : std_logic;
    signal l1_totem_2 : std_logic;
    signal l1_totem_4 : std_logic;
    signal l1_zdcm : std_logic;
    signal l1_zdcp : std_logic;
    signal l1_zdcm_bptx_and : std_logic;
    signal l1_zdcp_bptx_and : std_logic;
    signal l1_zdcm_zdcp_bptx_and : std_logic;
    signal l1_zdc_or_or_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_zdc_or_or_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_zdc_and_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_zdc_and_or_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_zdc_and_or_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_zdc_and_or_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_always_true : std_logic;
    signal l1_zero_bias : std_logic;
    signal l1_zero_bias_copy : std_logic;
    signal l1_bptx_or : std_logic;
    signal l1_not_bptx_or : std_logic;
    signal l1_isolated_bunch : std_logic;
    signal l1_first_bunch_in_train : std_logic;
    signal l1_second_bunch_in_train : std_logic;
    signal l1_last_bunch_in_train : std_logic;
    signal l1_first_bunch_after_train : std_logic;
    signal l1_first_bunch_before_train : std_logic;
    signal l1_second_last_bunch_in_train : std_logic;
    signal l1_first_collision_in_orbit : std_logic;
    signal l1_first_collision_in_orbit_centrality30_100_bptx_and : std_logic;
    signal l1_minimum_bias_hf0_and_bptx_and : std_logic;
    signal l1_not_minimum_bias_hf0_and_bptx_and : std_logic;
    signal l1_not_minimum_bias_hf0_or_bptx_and : std_logic;
    signal l1_minimum_bias_hf0_or_bptx_and : std_logic;
    signal l1_not_minimum_bias_hf0_and_bptx_and_totem_1 : std_logic;
    signal l1_not_minimum_bias_hf0_and_bptx_and_totem_2 : std_logic;
    signal l1_not_minimum_bias_hf0_and_bptx_and_totem_4 : std_logic;
    signal l1_not_minimum_bias_hf0_or_bptx_and_totem_1 : std_logic;
    signal l1_not_minimum_bias_hf0_or_bptx_and_totem_2 : std_logic;
    signal l1_not_minimum_bias_hf0_or_bptx_and_totem_4 : std_logic;
    signal l1_minimum_bias_hf1_and : std_logic;
    signal l1_minimum_bias_hf1_or : std_logic;
    signal l1_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_minimum_bias_hf1_xor_bptx_and : std_logic;
    signal l1_minimum_bias_hf1_and_or_ett10_bptx_and : std_logic;
    signal l1_not_minimum_bias_hf1_and : std_logic;
    signal l1_not_minimum_bias_hf1_or : std_logic;
    signal l1_not_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_minimum_bias_hf2_and : std_logic;
    signal l1_minimum_bias_hf2_or : std_logic;
    signal l1_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_not_minimum_bias_hf2_and : std_logic;
    signal l1_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_not_minimum_bias_hf2_or : std_logic;
    signal l1_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_centrality_30_100 : std_logic;
    signal l1_centrality_50_100 : std_logic;
    signal l1_centrality_20_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_centrality_30_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu_open_bptx_and : std_logic;
    signal l1_single_mu0_bptx_and : std_logic;
    signal l1_single_mu3_bptx_and : std_logic;
    signal l1_single_mu5_bptx_and : std_logic;
    signal l1_single_mu7_bptx_and : std_logic;
    signal l1_single_mu12_bptx_and : std_logic;
    signal l1_single_mu16_bptx_and : std_logic;
    signal l1_single_mu_open_centrality_70_100_bptx_and : std_logic;
    signal l1_single_mu3_centrality_70_100_bptx_and : std_logic;
    signal l1_single_mu_open_centrality_80_100_bptx_and : std_logic;
    signal l1_single_mu3_centrality_80_100_bptx_and : std_logic;
    signal l1_single_mu3_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu5_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu7_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu12_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu16_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu_open_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_mu0_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_mu3_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_mu_open_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_mu0_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_mu_open_centrality_70_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu_open_centrality_80_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet28_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet44_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet56_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu_open_single_jet64_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu3_single_jet28_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu3_single_jet32_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu3_single_jet40_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_mu3_single_eg12_bptx_and : std_logic;
    signal l1_single_mu_open_single_eg15_bptx_and : std_logic;
    signal l1_single_mu3_single_eg20_bptx_and : std_logic;
    signal l1_single_mu3_single_eg30_bptx_and : std_logic;
    signal l1_single_mu5_single_eg10_bptx_and : std_logic;
    signal l1_single_mu5_single_eg12_bptx_and : std_logic;
    signal l1_single_mu5_single_eg15_bptx_and : std_logic;
    signal l1_single_mu5_single_eg20_bptx_and : std_logic;
    signal l1_single_mu7_single_eg7_bptx_and : std_logic;
    signal l1_single_mu7_single_eg10_bptx_and : std_logic;
    signal l1_single_mu7_single_eg12_bptx_and : std_logic;
    signal l1_single_mu7_single_eg15_bptx_and : std_logic;
    signal l1_single_mu12_single_eg7_bptx_and : std_logic;
    signal l1_double_mu_open_bptx_and : std_logic;
    signal l1_double_mu_open_os_bptx_and : std_logic;
    signal l1_double_mu_open_ss_bptx_and : std_logic;
    signal l1_double_mu0_bptx_and : std_logic;
    signal l1_double_mu10_bptx_and : std_logic;
    signal l1_double_mu_open_max_dr2p0_bptx_and : std_logic;
    signal l1_double_mu_open_max_dr2p0_os_bptx_and : std_logic;
    signal l1_double_mu_open_max_dr3p5 : std_logic;
    signal l1_double_mu_open_max_dr3p5_bptx_and : std_logic;
    signal l1_double_mu0_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_double_mu_open_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_double_mu0_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_double_mu0_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_mu_open_centrality_10_100_bptx_and : std_logic;
    signal l1_double_mu_open_centrality_30_100_bptx_and : std_logic;
    signal l1_double_mu_open_centrality_40_100_bptx_and : std_logic;
    signal l1_double_mu_open_centrality_50_100_bptx_and : std_logic;
    signal l1_double_mu0_centrality_10_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_double_mu0_centrality_30_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_double_mu0_centrality_50_100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_single_jet8_bptx_and : std_logic;
    signal l1_single_jet16_bptx_and : std_logic;
    signal l1_single_jet24_bptx_and : std_logic;
    signal l1_single_jet28_bptx_and : std_logic;
    signal l1_single_jet32_bptx_and : std_logic;
    signal l1_single_jet36_bptx_and : std_logic;
    signal l1_single_jet40_bptx_and : std_logic;
    signal l1_single_jet44_bptx_and : std_logic;
    signal l1_single_jet48_bptx_and : std_logic;
    signal l1_single_jet56_bptx_and : std_logic;
    signal l1_single_jet60_bptx_and : std_logic;
    signal l1_single_jet64_bptx_and : std_logic;
    signal l1_single_jet72_bptx_and : std_logic;
    signal l1_single_jet80_bptx_and : std_logic;
    signal l1_single_jet8_fwd_bptx_and : std_logic;
    signal l1_single_jet16_fwd_bptx_and : std_logic;
    signal l1_single_jet28_fwd_bptx_and : std_logic;
    signal l1_single_jet36_fwd_bptx_and : std_logic;
    signal l1_single_jet44_fwd_bptx_and : std_logic;
    signal l1_single_jet56_fwd_bptx_and : std_logic;
    signal l1_single_jet64_fwd_bptx_and : std_logic;
    signal l1_single_jet8_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet16_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet24_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet28_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet32_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet36_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet40_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet44_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet48_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet56_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet60_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet64_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet8_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet16_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet24_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet28_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet32_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet36_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet40_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet44_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet48_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet56_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet60_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet64_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet8_fwd_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet16_fwd_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet28_fwd_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet36_fwd_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet44_fwd_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet56_fwd_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet64_fwd_centrality_30_100_bptx_and : std_logic;
    signal l1_single_jet8_fwd_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet16_fwd_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet28_fwd_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet36_fwd_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet44_fwd_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet56_fwd_centrality_50_100_bptx_and : std_logic;
    signal l1_single_jet64_fwd_centrality_50_100_bptx_and : std_logic;
    signal l1_double_jet16_and8_mid_eta2p7_bptx_and : std_logic;
    signal l1_double_jet16_and12_mid_eta2p7_bptx_and : std_logic;
    signal l1_double_jet20_and8_mid_eta2p7_bptx_and : std_logic;
    signal l1_double_jet20_and12_mid_eta2p7_bptx_and : std_logic;
    signal l1_double_jet28_and16_mid_eta2p7_bptx_and : std_logic;
    signal l1_double_jet16_and8_mid_eta2p7_centrality_30_100_bptx_and : std_logic;
    signal l1_double_jet16_and12_mid_eta2p7_centrality_30_100_bptx_and : std_logic;
    signal l1_double_jet20_and8_mid_eta2p7_centrality_30_100_bptx_and : std_logic;
    signal l1_double_jet20_and12_mid_eta2p7_centrality_30_100_bptx_and : std_logic;
    signal l1_double_jet28_and16_mid_eta2p7_centrality_30_100_bptx_and : std_logic;
    signal l1_double_jet16_and8_mid_eta2p7_centrality_50_100_bptx_and : std_logic;
    signal l1_double_jet16_and12_mid_eta2p7_centrality_50_100_bptx_and : std_logic;
    signal l1_double_jet20_and8_mid_eta2p7_centrality_50_100_bptx_and : std_logic;
    signal l1_double_jet20_and12_mid_eta2p7_centrality_50_100_bptx_and : std_logic;
    signal l1_double_jet28_and16_mid_eta2p7_centrality_50_100_bptx_and : std_logic;
    signal l1_single_eg3_bptx_and : std_logic;
    signal l1_single_eg5_bptx_and : std_logic;
    signal l1_single_eg7_bptx_and : std_logic;
    signal l1_single_eg12_bptx_and : std_logic;
    signal l1_single_eg15_bptx_and : std_logic;
    signal l1_single_eg21_bptx_and : std_logic;
    signal l1_single_eg30_bptx_and : std_logic;
    signal l1_single_iso_eg3_bptx_and : std_logic;
    signal l1_single_iso_eg7_bptx_and : std_logic;
    signal l1_single_iso_eg12_bptx_and : std_logic;
    signal l1_single_iso_eg15_bptx_and : std_logic;
    signal l1_single_iso_eg21_bptx_and : std_logic;
    signal l1_single_eg3_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_eg5_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_single_eg3_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_eg5_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_single_eg3_centrality_30_100_bptx_and : std_logic;
    signal l1_single_eg7_centrality_30_100_bptx_and : std_logic;
    signal l1_single_eg15_centrality_30_100_bptx_and : std_logic;
    signal l1_single_eg21_centrality_30_100_bptx_and : std_logic;
    signal l1_single_eg3_centrality_50_100_bptx_and : std_logic;
    signal l1_single_eg7_centrality_50_100_bptx_and : std_logic;
    signal l1_single_eg15_centrality_50_100_bptx_and : std_logic;
    signal l1_single_eg21_centrality_50_100_bptx_and : std_logic;
    signal l1_single_eg5_single_jet28_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg5_single_jet32_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg5_single_jet40_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg7_single_jet32_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg7_single_jet40_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg7_single_jet28_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg7_single_jet44_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg7_single_jet56_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg7_single_jet60_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg12_single_jet32_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg12_single_jet40_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg12_single_jet28_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg12_single_jet44_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg12_single_jet56_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg12_single_jet60_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg15_single_jet28_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg15_single_jet44_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg15_single_jet56_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg15_single_jet60_mid_eta2p7_bptx_and : std_logic;
    signal l1_single_eg15_single_jet28_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg15_single_jet44_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg15_single_jet56_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_single_eg15_single_jet60_mid_eta2p7_min_dr0p4_bptx_and : std_logic;
    signal l1_double_eg2_bptx_and : std_logic;
    signal l1_double_eg5_bptx_and : std_logic;
    signal l1_double_eg8_bptx_and : std_logic;
    signal l1_double_eg10_bptx_and : std_logic;
    signal l1_double_eg2_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_double_eg5_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_double_eg2_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_double_eg5_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_ett_asym40 : std_logic;
    signal l1_ett_asym50 : std_logic;
    signal l1_ett_asym60 : std_logic;
    signal l1_ett_asym70 : std_logic;
    signal l1_ett_asym80 : std_logic;
    signal l1_ett_asym40_bptx_and : std_logic;
    signal l1_ett_asym50_bptx_and : std_logic;
    signal l1_ett_asym60_bptx_and : std_logic;
    signal l1_ett_asym70_bptx_and : std_logic;
    signal l1_ett_asym80_bptx_and : std_logic;
    signal l1_ett_asym40_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett_asym50_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett_asym60_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett_asym70_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett_asym80_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett_asym40_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett_asym50_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett_asym60_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett_asym70_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett_asym80_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett5_bptx_and : std_logic;
    signal l1_ett5_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett5_not_minimum_bias_hf2_or : std_logic;
    signal l1_ett5_ett_asym40_bptx_and : std_logic;
    signal l1_ett5_ett_asym50_bptx_and : std_logic;
    signal l1_ett5_ett_asym60_bptx_and : std_logic;
    signal l1_ett5_ett_asym70_bptx_and : std_logic;
    signal l1_ett5_ett_asym80_bptx_and : std_logic;
    signal l1_ett5_ett_asym50_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett8_ett_asym50_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett8_ett_asym55_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett8_ett_asym60_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett8_ett_asym65_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett8_ett_asym70_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett8_ett_asym80_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett10_ett_asym50_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett10_ett_asym55_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym40_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym50_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym55_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym60_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym65_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym70_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym80_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym40_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym50_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym60_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym70_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett50_ett_asym80_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett60_ett_asym60_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett60_ett_asym65_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett65_ett_asym70_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett65_ett_asym80_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_ett5_not_ett30_bptx_and : std_logic;
    signal l1_ett35_not_ett80_bptx_and : std_logic;
    signal l1_ett40_not_ett95_bptx_and : std_logic;
    signal l1_ett45_not_ett110_bptx_and : std_logic;
    signal l1_ett50_not_ett120_bptx_and : std_logic;
    signal l1_ett55_not_ett130_bptx_and : std_logic;
    signal l1_not_ett20_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_not_ett80_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_not_ett95_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_not_ett20_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_not_ett80_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_not_ett95_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_not_ett20_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_not_ett80_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_not_ett95_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_not_ett100_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_not_ett150_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_not_ett200_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_not_ett110_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_not_ett110_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_not_ett150_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_not_ett150_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_castor_medium_jet : std_logic;
    signal l1_castor_medium_jet_bptx_and : std_logic;
    signal l1_castor_medium_jet_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_castor_medium_jet_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_castor_medium_jet_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_castor_medium_jet_single_mu0_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_castor_medium_jet_single_eg5_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_castor_muon : std_logic;
    signal l1_castor_muon_bptx_and : std_logic;
    signal l1_castor_high_jet : std_logic;
    signal l1_castor_high_jet_bptx_and : std_logic;
    signal l1_castor_high_jet_minimum_bias_hf1_or_bptx_and : std_logic;
    signal l1_castor_high_jet_not_minimum_bias_hf2_and_bptx_and : std_logic;
    signal l1_castor_high_jet_not_minimum_bias_hf2_or_bptx_and : std_logic;
    signal l1_castor_high_jet_or_minimum_bias_hf1_and_bptx_and : std_logic;
    signal l1_castor_high_jet_or_minimum_bias_hf2_and_bptx_and : std_logic;

-- ========================================================