-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2020_v0_1_8_massdr

-- Unique ID of L1 Trigger Menu:
-- 4df5c4be-8aa3-464e-a6b0-ea95c8c989e6

-- Unique ID of firmware implementation:
-- 575fd5ae-10e9-41f3-a476-6c3c08f40a9d

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.11.1

-- tmEventSetup version
-- v0.9.1

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        491, -- module_index: 0, name: L1_BPTX_BeamGas_B1_VME
        483, -- module_index: 1, name: L1_BPTX_OR_Ref3_VME
        479, -- module_index: 2, name: L1_FirstCollisionInTrain
        503, -- module_index: 3, name: L1_TOTEM_1
        469, -- module_index: 4, name: L1_UnpairedBunchBptxMinus
        426, -- module_index: 5, name: L1_ETMHF150
        260, -- module_index: 6, name: L1_ETT35
        400, -- module_index: 7, name: L1_HTT200er
          0, -- module_index: 8, name: L1_SingleMuCosmics
         19, -- module_index: 9, name: L1_SingleMu22
         11, -- module_index: 10, name: L1_SingleMu7_DQ
        174, -- module_index: 11, name: L1_SingleEG60
        314, -- module_index: 12, name: L1_SingleJet200
        311, -- module_index: 13, name: L1_SingleJet90
        305, -- module_index: 14, name: L1_Mu0upt100
        304, -- module_index: 15, name: L1_Mu0upt50
        157, -- module_index: 16, name: L1_Mu0upt20ip03
        155, -- module_index: 17, name: L1_Mu0upt20ip2
          1, -- module_index: 18, name: L1_SingleMuCosmics_BMTF
        306, -- module_index: 19, name: L1_SingleMuOpenupt5
         13, -- module_index: 20, name: L1_SingleMu12_DQ_BMTF
         32, -- module_index: 21, name: L1_SingleMu16er1p5
         25, -- module_index: 22, name: L1_SingleMu6er1p5
         28, -- module_index: 23, name: L1_SingleMu9er1p5
         41, -- module_index: 24, name: L1_DoubleMu0_SQ
        366, -- module_index: 25, name: L1_DoubleJet_80_30_Mass_Min420_DoubleMu0_SQ
        365, -- module_index: 26, name: L1_DoubleJet_80_30_Mass_Min420_Mu8
         89, -- module_index: 27, name: L1_QuadMu0
         90, -- module_index: 28, name: L1_QuadMu0_SQ
        109, -- module_index: 29, name: L1_DoubleMu4_SQ_EG9er2p5
        110, -- module_index: 30, name: L1_DoubleMu5_SQ_EG9er2p5
        205, -- module_index: 31, name: L1_DoubleEG_15_10_er2p5
        207, -- module_index: 32, name: L1_DoubleEG_22_10_er2p5
        209, -- module_index: 33, name: L1_DoubleEG_25_14_er2p5
        388, -- module_index: 34, name: L1_DoubleEG_5_er1p2
        390, -- module_index: 35, name: L1_DoubleEG_7_er1p2
        392, -- module_index: 36, name: L1_DoubleEG_9_er1p2
        342, -- module_index: 37, name: L1_DoubleJet120er2p5
        267, -- module_index: 38, name: L1_DoubleTau70er2p1
        327, -- module_index: 39, name: L1_SingleJet120_FWD3p0
        326, -- module_index: 40, name: L1_SingleJet90_FWD3p0
        214, -- module_index: 41, name: L1_DoubleEG_LooseIso22_12_er2p5
        269, -- module_index: 42, name: L1_DoubleIsoTau28er2p1
        271, -- module_index: 43, name: L1_DoubleIsoTau32er2p1
        273, -- module_index: 44, name: L1_DoubleIsoTau36er2p1
        218, -- module_index: 45, name: L1_DoubleLooseIsoEG24er2p1
        177, -- module_index: 46, name: L1_SingleLooseIsoEG28_FWD2p5
        224, -- module_index: 47, name: L1_TripleEG_16_12_8_er2p5
        226, -- module_index: 48, name: L1_TripleEG_18_17_8_er2p5
        374, -- module_index: 49, name: L1_TripleJet_105_85_75_DoubleJet_85_75_er2p5
        298, -- module_index: 50, name: L1_QuadJet36er2p5_IsoTau52er2p1
        346, -- module_index: 51, name: L1_DoubleJet112er2p3_dEta_Max1p6
         63, -- module_index: 52, name: L1_DoubleMu4p5_SQ_OS_dR_Max1p2
         58, -- module_index: 53, name: L1_DoubleMu0er1p5_SQ_OS_dR_Max1p4
         54, -- module_index: 54, name: L1_DoubleMu0er2p0_SQ_OS_dR_Max1p4
         50, -- module_index: 55, name: L1_DoubleMu_15_7_Mass_Min1
        433, -- module_index: 56, name: L1_DoubleEG_5_er1p2_dR_Max0p9
        121, -- module_index: 57, name: L1_Mu3_Jet16er2p5_dR_Max0p4
        135, -- module_index: 58, name: L1_Mu12er2p3_Jet40er2p3_dR_Max0p4_DoubleJet40er2p3_dEta_Max1p6
        143, -- module_index: 59, name: L1_DoubleMu3_dR_Max1p6_Jet90er2p5_dR_Max0p8
        274, -- module_index: 60, name: L1_DoubleIsoTau28er2p1_Mass_Max90
        236, -- module_index: 61, name: L1_LooseIsoEG30er2p1_Jet34er2p5_dR_Min0p3
    others => 0
);

-- ========================================================