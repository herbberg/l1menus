-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_Cidada_test_v1

-- Unique ID of L1 Trigger Menu:
-- 0cf00a60-7768-4152-bb84-6876899645a2

-- Unique ID of firmware implementation:
-- bdd2a2ac-dd4c-4029-a458-4a077c9988b5

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.15.0

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_jet_i3 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_jet60 : std_logic;

-- ========================================================