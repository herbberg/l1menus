-- ========================================================
-- from VHDL producer:

-- Module ID: 1

-- Name of L1 Trigger Menu:
-- L1Menu_adt_v4

-- Unique ID of L1 Trigger Menu:
-- 3ad635ba-a02d-467b-84ef-1022d6178c50

-- Unique ID of firmware implementation:
-- 842acd21-8068-4f00-a4d1-de71a487fb64

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.14.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i2 : std_logic;

-- Signal definition for algorithms names
    signal l1_adt_100 : std_logic;

-- ========================================================