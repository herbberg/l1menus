-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_simple_2

-- Unique ID of L1 Trigger Menu:
-- 4e10b5b5-9c10-4dbb-830e-c81310be9f45

-- Unique ID of firmware implementation:
-- 421b4fa7-8031-4747-b5fd-957f5dc307db

-- Scale set:
-- scales_2024_05_15

-- VHDL producer
-- version: 2.20.1
-- hash value: 37aeed0f04da76b667e2567c8eee7fb6e0bbfdcc7e4a47a65d22d7168cf55357

-- tmEventSetup
-- version: 0.13.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_htt_i3 : std_logic;

-- Signal definition for algorithms names
    signal l1_htt120er : std_logic;

-- ========================================================