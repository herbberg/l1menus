-- ========================================================
-- from VHDL producer:

-- Module ID: 2

-- Name of L1 Trigger Menu:
-- L1Menu_Cidada_test_v2

-- Unique ID of L1 Trigger Menu:
-- ded9c4b7-1624-4694-93ed-c9e7bf41a550

-- Unique ID of firmware implementation:
-- a6af76db-ec42-4888-8409-d2323ca95556

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.15.0

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_eg_i0 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_eg3 : std_logic;

-- ========================================================