-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2022_adt_test

-- Unique ID of L1 Trigger Menu:
-- 9f50db6e-c51d-40e2-8252-459006e512fc

-- Unique ID of firmware implementation:
-- 7d77f46e-1e11-4138-b324-80855db4e2e1

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.12.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- -- Signal definition for conditions names
--     signal single_mu_i0 : std_logic;
--
-- -- Signal definition for algorithms names
--     signal l1_single_mu0 : std_logic;

-- Signal definition for conditions names
    signal adt_sig : std_logic;

-- Signal definition for algorithms names
    signal l1_adt : std_logic;

-- ========================================================
