-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_Collisions2022_adt_test_ext_sig_v2

-- Unique ID of L1 Trigger Menu:
-- b581e141-1a2d-45fa-81d7-45348fab94a3

-- Unique ID of firmware implementation:
-- e8c3c770-2d65-44e6-bcd7-da256a4cb74f

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.14.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i5 : std_logic;

-- Signal definition for algorithms names
    signal l1_adt_5 : std_logic;

-- ========================================================