-- ========================================================
-- from VHDL producer:

-- Module ID: 5

-- Name of L1 Trigger Menu:
-- L1Menu_Cicada_Adt_Topo_test

-- Unique ID of L1 Trigger Menu:
-- e50b8093-a248-4fd5-baf6-5b197178654a

-- Unique ID of firmware implementation:
-- 7fe6a178-b7c7-4223-a477-aecdf8df542c

-- Scale set:
-- scales_2024_01_04

-- VHDL producer version
-- v2.17.0

-- tmEventSetup version
-- v0.12.0

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
         10, -- module_index: 0, name: L1_TOPO_1006_ext
          3, -- module_index: 1, name: L1_CICADA_10p023
          2, -- module_index: 2, name: L1_CICADA_142p273
    others => 0
);

-- ========================================================