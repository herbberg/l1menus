-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_calo_comp_pt_obj_nr_condition_test_v2

-- Unique ID of L1 Trigger Menu:
-- f9f63b7d-bf5d-4d02-a79c-e1a228890ebe

-- Unique ID of firmware implementation:
-- ffa7fad4-8dd6-4707-a137-cceafccc2fe0

-- Scale set:
-- scales_2024_02_14

-- VHDL producer
-- version: 2.18.0
-- hash value: 1c5712f4e1570ec4dd437d604d3d1604f5a84fd8a70cb4ddfc66cba619604f7a

-- tmEventSetup
-- version: 0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    --signal quad_jet_i5 : std_logic;
    signal six_jets_i1 : std_logic;

-- Signal definition for algorithms names
    signal l1_six_jets_23 : std_logic;

-- ========================================================
