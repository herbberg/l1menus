-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_Cicada_Adt_Topo_test

-- Unique ID of L1 Trigger Menu:
-- e50b8093-a248-4fd5-baf6-5b197178654a

-- Unique ID of firmware implementation:
-- 7fe6a178-b7c7-4223-a477-aecdf8df542c

-- Scale set:
-- scales_2024_01_04

-- VHDL producer version
-- v2.17.0

-- tmEventSetup version
-- v0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal anomaly_detection_trigger_i10 : std_logic;
    signal single_eg_i6 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_eg8er2p5 : std_logic;
    signal l1_adt_174 : std_logic;

-- ========================================================