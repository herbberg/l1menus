-- ========================================================
-- from VHDL producer:

-- Module ID: 2

-- Name of L1 Trigger Menu:
-- L1Menu_test_esums_instances_v1

-- Unique ID of L1 Trigger Menu:
-- f7b5ee69-e72e-4011-aa54-9fdcb44159a6

-- Unique ID of firmware implementation:
-- 6f3e759e-dcce-42f7-afca-398c7df773ad

-- Scale set:
-- scales_2017_05_23

-- VHDL producer version
-- v2.7.3

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
        421, -- module_index: 0, name: L1_ETMHF100
        444, -- module_index: 1, name: L1_ETMHF110_HTT60er_NotSecondBunchInTrain
        461, -- module_index: 2, name: L1_MinimumBiasHF0_AND_BptxAND
        150, -- module_index: 3, name: L1_DoubleMu3_SQ_HTT220er
        151, -- module_index: 4, name: L1_DoubleMu3_SQ_HTT240er
        428, -- module_index: 5, name: L1_ETMHF90_HTT60er
        152, -- module_index: 6, name: L1_DoubleMu3_SQ_HTT260er
        145, -- module_index: 7, name: L1_DoubleMu3_SQ_ETMHF50_HTT60er
        132, -- module_index: 8, name: L1_Mu6_HTT250er
        424, -- module_index: 9, name: L1_ETMHF130
        148, -- module_index: 10, name: L1_DoubleMu3_SQ_ETMHF60_Jet60er2p5
        432, -- module_index: 11, name: L1_ETMHF130_HTT60er
        422, -- module_index: 12, name: L1_ETMHF110
        423, -- module_index: 13, name: L1_ETMHF120
        443, -- module_index: 14, name: L1_ETMHF120_NotSecondBunchInTrain
        430, -- module_index: 15, name: L1_ETMHF110_HTT60er
        146, -- module_index: 16, name: L1_DoubleMu3_SQ_ETMHF50_Jet60er2p5_OR_DoubleJet40er2p5
        131, -- module_index: 17, name: L1_Mu6_HTT240er
        147, -- module_index: 18, name: L1_DoubleMu3_SQ_ETMHF50_Jet60er2p5
        431, -- module_index: 19, name: L1_ETMHF120_HTT60er
        429, -- module_index: 20, name: L1_ETMHF100_HTT60er
    others => 0
);

-- ========================================================