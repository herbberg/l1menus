-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_1_0_utm_0_11_zdc

-- Unique ID of L1 Trigger Menu:
-- c1d5a598-16e4-45bf-8da2-398033004599

-- Unique ID of firmware implementation:
-- 57c2bcc2-8b13-46b5-b0fc-8673f5867e06

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.1

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i3 : std_logic;
    signal single_ext_i34 : std_logic;
    signal single_ext_i79 : std_logic;
    signal single_ext_i8 : std_logic;
    signal single_htt_i36 : std_logic;
    signal single_eg_i52 : std_logic;
    signal single_jet_i65 : std_logic;
    signal single_mu_i69 : std_logic;
    signal single_mu_i71 : std_logic;
    signal single_mu_i76 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_and_ref4_vme : std_logic;
    signal l1_bptx_not_or_vme : std_logic;
    signal l1_first_collision_in_train : std_logic;
    signal l1_htt200er : std_logic;
    signal l1_single_eg10er2p5 : std_logic;
    signal l1_single_jet35er2p5 : std_logic;
    signal l1_single_mu0_dq : std_logic;
    signal l1_single_mu0_omtf : std_logic;
    signal l1_single_mu_cosmics_bmtf : std_logic;
    signal l1_unpaired_bunch_bptx_minus : std_logic;

-- ========================================================