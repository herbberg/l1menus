-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2018_v4_2_0_new_scale

-- Unique ID of L1 Trigger Menu:
-- 786b195b-7fe4-4c23-a571-ac5068c6fa09

-- Unique ID of firmware implementation:
-- 16aa0ff4-bb99-4e7c-93a6-91d053a5e21c

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.12.1

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i197 : std_logic;
    signal single_ext_i59 : std_logic;
    signal single_ext_i86 : std_logic;
    signal single_ext_i92 : std_logic;
    signal single_ett_i55 : std_logic;
    signal single_htt_i53 : std_logic;
    signal single_eg_i28 : std_logic;
    signal single_eg_i30 : std_logic;
    signal single_jet_i41 : std_logic;
    signal single_jet_i46 : std_logic;
    signal single_jet_i47 : std_logic;
    signal single_mu_i1 : std_logic;
    signal single_mu_i8 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_mu_cosmics_bmtf : std_logic;
    signal l1_single_mu0_omtf : std_logic;
    signal l1_single_eg50 : std_logic;
    signal l1_single_eg10er2p5 : std_logic;
    signal l1_single_jet35er2p5 : std_logic;
    signal l1_single_jet60_fwd3p0 : std_logic;
    signal l1_htt360er : std_logic;
    signal l1_ett2000 : std_logic;
    signal l1_totem_3 : std_logic;
    signal l1_bptx_not_or_vme : std_logic;
    signal l1_bptx_and_ref4_vme : std_logic;
    signal l1_castor1 : std_logic;

-- ========================================================