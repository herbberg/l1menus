-- ========================================================
-- from VHDL producer:

-- Module ID: 3

-- Name of L1 Trigger Menu:
-- L1Menu_adt_v7

-- Unique ID of L1 Trigger Menu:
-- 63d8f700-507a-4a7b-bde4-58b4c3437959

-- Unique ID of firmware implementation:
-- ff999d54-d3e2-4483-8c05-b631978b815b

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.14.0

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i7 : std_logic;

-- Signal definition for algorithms names
    signal l1_adt_80 : std_logic;

-- ========================================================