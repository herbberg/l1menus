-- ========================================================
-- from VHDL producer:

-- Module ID: 1

-- Name of L1 Trigger Menu:
-- L1Menu_calo_comp_pt_obj_nr_condition_test

-- Unique ID of L1 Trigger Menu:
-- b64d6c4c-db5f-46a5-b59c-3159102b5b6d

-- Unique ID of firmware implementation:
-- cd5c3e0b-538f-44eb-aa06-4ee14281d9ca

-- Scale set:
-- scales_2024_02_14

-- VHDL producer
-- version: 2.18.0
-- hash value: 1c5712f4e1570ec4dd437d604d3d1604f5a84fd8a70cb4ddfc66cba619604f7a

-- tmEventSetup
-- version: 0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_eg_i1 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_eg10er2p5 : std_logic;

-- ========================================================