-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_utm_0_11_test_v3

-- Unique ID of L1 Trigger Menu:
-- 36a2b4c9-da1a-4698-be00-93a32f4e85dc

-- Unique ID of firmware implementation:
-- d3f20e01-a22f-46d2-b314-c95247e5ac55

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.0

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i2 : std_logic;
    signal zdc_plus_i11 : std_logic;

-- Signal definition for algorithms names
    signal l1_adt_4000_ext : std_logic;
    signal l1_zdc_plus_128 : std_logic;

-- ========================================================