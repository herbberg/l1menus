-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_test_orm

-- Unique ID of L1 Trigger Menu:
-- 6b3c4161-f14b-4d94-abd9-6ac0308248ac

-- Unique ID of firmware implementation:
-- d0109e5f-d8d0-4715-8a9c-0fd5e15f0dd5

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.11.1

-- tmEventSetup version
-- v0.9.1

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
          0, -- module_index: 0, name: L1_DoubleJet35_Dphi_0_1_IsoTau45_RmOvlp
    others => 0
);

-- ========================================================