-- ========================================================
-- from VHDL producer:

-- Module ID: 2

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2022_v1_1_0_utm_0_11_zdc

-- Unique ID of L1 Trigger Menu:
-- e3e2c317-bee5-4ffa-8bd7-765abf589aa1

-- Unique ID of firmware implementation:
-- b54ce0e7-99c8-4d78-ace7-3e12ebd64fc5

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.1

-- tmEventSetup version
-- v0.11.2

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_ext_i10 : std_logic;
    signal single_ext_i5 : std_logic;
    signal muon_shower0_i16 : std_logic;
    signal single_htt_i38 : std_logic;
    signal single_eg_i56 : std_logic;
    signal single_jet_i57 : std_logic;
    signal single_jet_i63 : std_logic;
    signal single_jet_i64 : std_logic;
    signal single_mu_i68 : std_logic;
    signal single_mu_i72 : std_logic;

-- Signal definition for algorithms names
    signal l1_bptx_beam_gas_b2_vme : std_logic;
    signal l1_bptx_or_ref4_vme : std_logic;
    signal l1_mu_shower_one_nominal : std_logic;
    signal l1_htt360er : std_logic;
    signal l1_single_eg8er2p5 : std_logic;
    signal l1_single_jet120 : std_logic;
    signal l1_single_jet35_fwd3p0 : std_logic;
    signal l1_single_mu0_bmtf : std_logic;
    signal l1_single_mu22 : std_logic;

-- ========================================================