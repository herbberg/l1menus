-- ========================================================
-- from VHDL producer:

-- Module ID: 1

-- Name of L1 Trigger Menu:
-- L1Menu_Cicada_test_16bits_v2

-- Unique ID of L1 Trigger Menu:
-- e50b8093-a248-4fd5-baf6-5b197178654a

-- Unique ID of firmware implementation:
-- 62d16def-def4-49df-a36a-08b0f2187b5f

-- Scale set:
-- scales_2023_12_14

-- VHDL producer version
-- v2.17.0

-- tmEventSetup version
-- v0.12.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_eg_i6 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_eg8er2p5 : std_logic;

-- ========================================================