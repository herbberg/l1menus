-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_CollisionsHeavyIons2018_v4_2_0_new_scale

-- Unique ID of L1 Trigger Menu:
-- 786b195b-7fe4-4c23-a571-ac5068c6fa09

-- Unique ID of firmware implementation:
-- 16aa0ff4-bb99-4e7c-93a6-91d053a5e21c

-- Scale set:
-- scales_2021_03_02

-- VHDL producer version
-- v2.12.1

-- tmEventSetup version
-- v0.10.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal single_cent7_i99 : std_logic;
    signal single_ext_i69 : std_logic;
    signal single_ext_i87 : std_logic;
    signal single_ext_i95 : std_logic;
    signal single_htt_i50 : std_logic;
    signal single_eg_i31 : std_logic;
    signal single_jet_i39 : std_logic;
    signal single_jet_i43 : std_logic;
    signal single_mu_i0 : std_logic;
    signal single_mu_i19 : std_logic;
    signal single_mu_i7 : std_logic;

-- Signal definition for algorithms names
    signal l1_single_mu_cosmics : std_logic;
    signal l1_single_mu0_bmtf : std_logic;
    signal l1_single_mu22_emtf : std_logic;
    signal l1_single_eg15er2p5 : std_logic;
    signal l1_single_jet120 : std_logic;
    signal l1_single_jet60er2p5 : std_logic;
    signal l1_htt120er : std_logic;
    signal l1_unpaired_bunch_bptx_minus : std_logic;
    signal l1_bptx_or_ref3_vme : std_logic;
    signal l1_bptx_beam_gas_b1_vme : std_logic;
    signal l1_centrality_saturation : std_logic;

-- ========================================================