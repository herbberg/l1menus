-- ========================================================
-- from VHDL producer:

-- Module ID: 0

-- Name of L1 Trigger Menu:
-- L1Menu_test_invmass_div_dr

-- Unique ID of L1 Trigger Menu:
-- 3c0c7341-bcb2-4f71-9732-a11cb177c360

-- Unique ID of firmware implementation:
-- 9b489ec0-fbf4-4941-985c-52e06058d80c

-- Scale set:
-- scales_2018_08_07

-- VHDL producer version
-- v2.8.0

-- ********************************************************************
-- Created manually for muon_muon_corr_cond (mass_div_dr) and calo_calo_corr_cond
-- ********************************************************************

-- HB 2016-09-16: constants for algo_mapping_rop.
type global_index_array is array (0 to NR_ALGOS-1) of integer;
constant global_index: global_index_array := (
          0, -- module_index: 0, name: l1_muon_invmass_div_dr_1
          1, -- module_index: 1, name: l1_muon_invmass_div_dr_2
          2, -- module_index: 2, name: l1_double_jet30er2p5_mass_min330_d_eta_max1p5
          3, -- module_index: 3, name: l1_double_jet45_mass_min620
    others => 0
);

-- ========================================================
