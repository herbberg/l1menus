-- ========================================================
-- from VHDL producer:

-- Module ID: 4

-- Name of L1 Trigger Menu:
-- L1Menu_utm_0_11_test

-- Unique ID of L1 Trigger Menu:
-- 36a2b4c9-da1a-4698-be00-93a32f4e85dc

-- Unique ID of firmware implementation:
-- e605ff0a-13b6-419c-891b-16096a11f0b8

-- Scale set:
-- scales_2023_02_16

-- VHDL producer version
-- v2.14.0

-- tmEventSetup version
-- v0.11.0

-- Signal definition of pt, eta and phi for correlation conditions.

-- Signal definition for cuts of correlation conditions.

-- Signal definition for muon charge correlations.

-- Signal definition for conditions names
    signal zdc_minus_i7 : std_logic;
    signal single_mu_i4 : std_logic;

-- Signal definition for algorithms names
    signal l1_zdc_minus_60 : std_logic;
    signal l1_single_mu_index_4_8 : std_logic;

-- ========================================================